/*module oscill_sim(level, sample, slope, mode, rst, clk, trig_en, asghar, norm_trig);
input unsigned [7:0] level, sample;
input slope, mode, rst, clk;
output trig_en, norm_trig;
output [19:0] asghar;
trig tr(level, sample, slope, mode, rst, clk, trig_en, asghar, norm_trig);
endmodule*/

module oscill_sim();
endmodule